end gr_controller;
