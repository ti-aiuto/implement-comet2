library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity prom is
	port(
		P_COUNT : in std_logic_vector(15 downto 0);
		PROM_OUT : out std_logic_vector(15 downto 0)
	);
end prom;

architecture RTL of prom is

subtype WORD is std_logic_vector(0 to 15);

type MEMORY is array (0 to 31) of WORD;

constant MEM : MEMORY := 
	(
		"0001001000010000", -- LAD GR1 64
		"0000000001000000", 
		"0001001000100000", -- LAD GR2 24
		"0000000000011000", 
		"0001010000110001", -- LD GR3 GR1
		"0001010001000010", -- LD GR4 GR2
		"0001010000010011", -- LD GR1 GR3 [LOOP1]
		"0001010000100100", -- LD GR2 GR4
		"0100010000010010", -- CPA GR1 GR2 [LOOP2]
		"0110001100000000", -- JZE OWARI
		"0000000000010100", 
		"0110000100000000", -- JMI NEXT
		"0000000000010000", 
		"0010010100010010", -- SUBA GR1 GR2
		"0110010000000000", -- JUMP LOOP2
		"0000000000001000", 
		"0001010000110010", -- LD GR3 GR2 [NEXT]
		"0001010001000001", -- LD GR4 GR1
		"0110010000000000", -- JUMP LOOP1
		"0000000000000110",
		"0001010000010010", -- LD GR1 GR2 [OWARI]
		"0000000000000000", -- NOP 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000"
	);

begin 
	PROM_OUT <= MEM(conv_integer(P_COUNT(4 downto 0)));
end RTL;
